====================================================================================================
No referer found for: sv domains
Tested domain: ayudaenaccion.org.sv
====================================================================================================
