====================================================================================================
No referer found for: sv domains
Tested domain: ayudaenaccion.org.sv
====================================================================================================
====================================================================================================
No referer found for: sv domains
Tested domain: upisss.gob.sv
====================================================================================================
